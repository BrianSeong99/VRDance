PK   ,d�V�hCwD  ��    cirkitFile.json��M�י�����J�{��zY��E�,3�(�j�"�n
T�/c��O��V�����,���?O���:?o���O�û��4|�~:_7o������z���˟�������2|{=~��y����O?}<���z:�s�̰{�^�^_�<����~�=�|}|��}{�o�~|��U�m�~���?���
�F�!�Іm�!�І]�!�І}�!�ІC�!�І�4CV���Y�6�N3d��&͐U5�A��E@T泲��2-1���2-1��3-1��#3-1��C3-1��c3-1��3-1��3-1���ggZb��ggZb� o4�ٹ�ggZb��ggZb��ggZb��ggZb��ggZb��ggZb��ggZb���LK���LK���LK����s��δ�H��δ�H��δ�H��δ�H��δ�H��δD���LK���LK���LK���LK��C�|v��ٙ�)�ٙ�)�ٙ�)�ٙ�)�ٙ�h�!��i��"��i��"��i��"��i��"��i��|E���C>;�#E>;�#E>;�#E>;�m��ggZb��ggZb��g�J�������x~��O9/������r��o�r��uK7	R����uK׆��nk��t�ҵag��Y�(]�tc����w��[��=���`��t�ҍ�oo����Q�n����z��zG麥k�k��k��떮o�wo�w��[��T ~s�����o:ψ���B��/:.7��1�t���[���o:����M��u�7�����a�:�Nc�p�|�Mg���uX����S��?�<,_�|��t�n��c��d=�����1�t' ������o�̀���p�8p���������u�7� ����a�:��`�p��|�M�v��X�����F�?�?,_�|�M)����c������1�t;�����u�7ݫ����a�:�nb�p��|�Mw����>f��������c���(����1�t�������o��������u�7�6����a�:��Ic�p��|�M7��{�?,_�|��t����c��V=����1��< ����c��I�?}�C_���c������1�������c���?�?,_�|�;��X����g�`�p��|�MOI��p��|�M�w����a�:曞L������u�7=S������oz����1��#쟾m�����q�������ozv����1���+����c��y]�?�?,_�|ӓƬw�X����g�a�p��|�MOw����a�z���Mp��{wy�\�s|�k��6/��PWBm��3DH�6�g���m��!�ی�!BB�Q?C��n�	�����"$t4DH��v�PD��v��r���VJ� ��Xvw�J������\)��r bb�Y�+�v[DL,Ƿ,Ǖ�<Z����o������R����-�q�4O"&��[��Ji�EDL,Ƿ,Ǖ�<���8���q�4�)"&�I��(�����R�����q�4�2"&��;��JilDL,��,Ǖ�<战X��Y�+�y�1���݇�,��,Ǖ�<	��X��Y�+�y.1�߳WJ�$������R�g&���q�4OP"&���z�����R��*���q�4Y"&��w,Ǖ�<r��X�߱�=�?~���9<�z;%T�s�\��N��>?�g�`]/f������
����q��}"�
}�`]/m��3���
��
�q���#�
}�`]/t��K���
��z�q��}%�
}�`]/{��c���
���q���&�
}�`]/��w�5�k������T�ڶ����ۢ�UӻV��^Vz[S�Jh�z���Jok�W	m[}zY�mM+�m�P/+���a%�m=�e��5U�����C�������ж�������T�ڶ���ۚZVB�zY��BM/+��T��������C�^Vz[��XM/[��zY�mM/+�Z���������^Vz[��Jh�aW/+���e%��諗������`��JokzY	m0�e��5���6����dRM/+�Ff���������^Vz[��Jh�qZ/+�-:�X��Vð^Vz[��Jh�Q[/+���e%��ୗ������`��JokzY	m0��e��5���6����ۚ^VB�zYy�������^Vz[��Jh�a^/+���e%��h��������`���Jo������՘��������`��JokzY	m0�e��5���6���ۚ^VB�{Y�mM/+������]��Jh�Qb/+���e%��`��������`���JokzY	m0t�e��5���6A���ۢ�|���� ��������`<��JokzY	m0��e��5���6]���ۚ^VB2{Y�d��^VB�5{Y�mM/+����������>�o#ϟ��O'0��x��t=>|	��F��P�m3"$4�<"$4�<"$4�<"$4�<"$4�<"$4�<"$4�<"$4�<"$��if�.�]l���,��R�������[)�y��0���,��R������B\)�y��0�߲WJ�ȳar��p��[��Jiy6L,Ƿ,Ǖ�2�l�X�oY�+�e��0�߲WJ�ȳ��,�w,Ǖ�2�l��')���;��Jiy6L,�w,Ǖ�2�l�X��X�+�e��0�߳WJ�ȳab9�g9����g��>w��߳WJ�ȳab9�g9����g��r|�r\)-#������Jiy6L,�,Ǖ�2�l�ܷ���M����Jiy6L,�,Ǖ�2�l�X�߱WJ�ȳab9~�r�����i��i>�:���ȳVe��n����|ā
�`�8�:ŧU�����3q`u�J�B_+X��g���V�V��V�#�āՍ*�
}�`F����TZ�Z��<V7��*���5y&�nQiU�kk0�LXݠҪ��
�`�ټ��)\��d���r�ж`6��Jo�jWM�Z�&sY�mM�*�m�l2����ԯ��&sY�mM+�m�l2����԰��&sY�mM+�m�l2����Ա��&sY�mM%+�m�l2����Բ�h���ojzY	m4��e��5���6y��ۢ��jz�z6��JokzY	m4��e��5���6y��ۚ^VB�<sY�mM/+��F���������F#�\Vz[��Jh��g.+���e%���3��'�jzY	m4��e��5���6y��ۚ^VB�<sY�m�qŚ^��M��ۚ^VB�<sY�mM/+��F���������F#�\Vz[��Jh��g.+���e%���3�������h��ʛ5���6y��ۚ^VB�<sY�mM/+��F���������F#�\Vz[t�����g���������F#�\Vz[��Jh��g.+���e%���3�������h��JokzY	m4��e���^VB�<sY�mM/+��F���������F#�\Vz[��Jh��g.+���e%���3���=棦��g���������F#�\Vz[��Jh��g.+���e%���3�������h���'+����h��JokzY	m4��e��5���iy1����w���u8���y�^l~8_O����w����8\������W_��ߺ���|?����}�ێ�����_���������L�ҟ��`Uz�қ?�'��h��$EZb^�NR�%���$EZb^�NR�%�e�$EZb^�NR�%��$EZb^}NR�%��$EZ�͛����)��g��h��r�dh!��h�r��hA��h�~r�dia��h�Nr����i^cYV�r����)��-�ӼƲ��� y�y��X֑� O� O��
r����i^cY;�VI��;��y�e�8�!��� Ow O��bq����i^cY&�r�<݁<�k,�Y��{��y�ei8��t�4��,
g9�g��CS��{��y�e-8��t�4���g9@��A��5������ O O���o����i^cY��r�o���P O O��Ro����i^cY��r�<�y��X�w� O�@��5��Q��Q*�7�EI���N�M�ֿ�9���|�nn����D9=���q��wu���,_���|��+'N��g������]]+qz�?���&_����#�Y�`�6�zW�C����;��׻����/أM���5�G��|��l���. ����;^]A0a�Z�����C֛�P�x��&l��*4�:�	[��
����`�l�BA㡮%����P�x��	&l�6*4�z�	[��
����`�l�BA㡮)�0Z`���j�S0a��
����`�hQ
�W&����H���P�L-�BA��)�0ZB���C�S0a�x
����`�h�
uO��т)4Ꞃ	��R(h<�=F��PМ�=FˣP�x�{
&�F���P�L-�BA�!?ޥ{�z�
uO���2(4Ꞃ	�P(h<�=FK�P�x�{
&�=���P�L-wBA��)�0Z脂���)�0Zℂ�C�S0a��	����`�hY
uO��т&4�(����'���P�L-bBA��)�0Z����C�S0a�p	����`�h�
uO���b%47uO���2%4Ꞃ	�J(h<�=FK�P�x�{
&�%���P�L-GBA�!�6�{�zs
uO���$4Ꞃ	��G(h<�=FˎP�x�{
&���y���)�0Zj���C�S0a������D���ؼ�|���xz|�����O�a?��������4�8L�����il|8~sz����a��р�������i��_m�%��ݰ����4��nx8��|�bS ����ǧ���������7O���3�޿����۟{�y���g?��>�?|���gN�o?L�s�~�����O��>�|��t��__�߯������|����˅�����=>������?�����t���O�=>~>>����>�����S�_�PK   ,d�V�hCwD  ��            ��    cirkitFile.jsonPK      =   q    